module fetch(input clock,
		input reset,
		input [3:0] state,
		input [15:0] taddr,
		input br_taken,
		output [15:0] pc,
		output [15:0] npc,
		output [15:0] rd);
endmodule